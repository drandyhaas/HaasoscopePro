// remoteupdate.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module remoteupdate (
		output wire        busy,        //        busy.busy
		input  wire        clock,       //       clock.clk
		output wire [28:0] data_out,    //    data_out.data_out
		input  wire [2:0]  param,       //       param.param
		input  wire        read_param,  //  read_param.read_param
		input  wire [1:0]  read_source, // read_source.read_source
		input  wire        reconfig,    //    reconfig.reconfig
		input  wire        reset,       //       reset.reset
		input  wire        reset_timer  // reset_timer.reset_timer
	);

	remoteupdate_remote_update_0 remote_update_0 (
		.busy        (busy),        //        busy.busy
		.data_out    (data_out),    //    data_out.data_out
		.param       (param),       //       param.param
		.read_param  (read_param),  //  read_param.read_param
		.reconfig    (reconfig),    //    reconfig.reconfig
		.reset_timer (reset_timer), // reset_timer.reset_timer
		.read_source (read_source), // read_source.read_source
		.clock       (clock),       //       clock.clk
		.reset       (reset)        //       reset.reset
	);

endmodule
