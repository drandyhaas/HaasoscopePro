// asmi.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module asmi (
		input  wire [23:0] addr,          //          addr.addr
		input  wire        bulk_erase,    //    bulk_erase.bulk_erase
		output wire        busy,          //          busy.busy
		input  wire        clkin,         //         clkin.clk
		output wire        data_valid,    //    data_valid.data_valid
		input  wire [7:0]  datain,        //        datain.datain
		output wire [7:0]  dataout,       //       dataout.dataout
		output wire        illegal_erase, // illegal_erase.illegal_erase
		output wire        illegal_write, // illegal_write.illegal_write
		input  wire        rden,          //          rden.rden
		input  wire        read,          //          read.read
		input  wire        reset,         //         reset.reset
		input  wire        write          //         write.write
	);

	asmi_asmi_parallel_0 asmi_parallel_0 (
		.clkin         (clkin),         //         clkin.clk
		.read          (read),          //          read.read
		.rden          (rden),          //          rden.rden
		.addr          (addr),          //          addr.addr
		.write         (write),         //         write.write
		.datain        (datain),        //        datain.datain
		.bulk_erase    (bulk_erase),    //    bulk_erase.bulk_erase
		.reset         (reset),         //         reset.reset
		.dataout       (dataout),       //       dataout.dataout
		.busy          (busy),          //          busy.busy
		.data_valid    (data_valid),    //    data_valid.data_valid
		.illegal_write (illegal_write), // illegal_write.illegal_write
		.illegal_erase (illegal_erase)  // illegal_erase.illegal_erase
	);

endmodule
